-- DECODER_PARALLEL
LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY simpleLogic;
USE simpleLogic.all;

ENTITY decoder_parallel IS
	PORT(